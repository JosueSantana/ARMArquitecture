module test_mux_16x1;
	wire [31:0] Y;
	reg [3:0] S;
	reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15;

	parameter sim_time = 200;
	mux_16x1 mux16(Y,S,I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15);
	initial #sim_time $finish;

	initial begin
		S = 4'b0000;
		I0 = 32'b00000000000000000000000000000000;
		I1 = 32'b00000000000000000000000000000001;
		I2 = 32'b00000000000000000000000000000010;
		I3 = 32'b00000000000000000000000000000011;
		I4 = 32'b00000000000000000000000000000100;
		I5 = 32'b00000000000000000000000000000101;
		I6 = 32'b00000000000000000000000000000110;
		I7 = 32'b00000000000000000000000000000111;
		I8 = 32'b00000000000000000000000000001000;
		I9 = 32'b00000000000000000000000000001001;
		I10= 32'b00000000000000000000000000001010;
		I11= 32'b00000000000000000000000000001011;
		I12= 32'b00000000000000000000000000001100;
		I13= 32'b00000000000000000000000000001101;
		I14= 32'b00000000000000000000000000001110;
		I15= 32'b00000000000000000000000000001111;

		repeat(16) #10 S=S+4'b0001;
	end

	initial begin
		$display(" S I0 I1 I2 I3 I4 I5 I6 I7 I8 I9 I10 I11 I12 I13 I14 I15 Y");
		$monitor(" %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b", S, I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, Y);
	end
endmodule
		