module control_unit (output reg regClr, marEn, irEn, memEn, memRW, input [31:0] status_reg, instruction, input [3:0] cond, input clr, clk);
	


endmodule